module main (
    input clk,
    input rst,
    input [7:0] phase, 
    input [31:0] desired_freq,   
    output reg signed [7:0] out 
);
parameter CLOCK_FREQUENCY = 100_000_000;

reg [7:0] phase_acc = 0; 
reg signed [7:0] lut [0:255];
reg [31:0] phase_increment; 

initial begin
    $readmemb("I:/FPGA/Vivado/dds_signed/main/main.srcs/sources_1/new/lut_values.txt", lut);
    /*
     lut[0] = 0;
lut[1] = 3;
lut[2] = 6;
lut[3] = 9;
lut[4] = 12;
lut[5] = 16;
lut[6] = 19;
lut[7] = 22;
lut[8] = 25;
lut[9] = 28;
lut[10] = 31;
lut[11] = 34;
lut[12] = 37;
lut[13] = 40;
lut[14] = 43;
lut[15] = 46;
lut[16] = 49;
lut[17] = 51;
lut[18] = 54;
lut[19] = 57;
lut[20] = 60;
lut[21] = 63;
lut[22] = 65;
lut[23] = 68;
lut[24] = 71;
lut[25] = 73;
lut[26] = 76;
lut[27] = 78;
lut[28] = 81;
lut[29] = 83;
lut[30] = 85;
lut[31] = 88;
lut[32] = 90;
lut[33] = 92;
lut[34] = 94;
lut[35] = 96;
lut[36] = 98;
lut[37] = 100;
lut[38] = 102;
lut[39] = 104;
lut[40] = 106;
lut[41] = 107;
lut[42] = 109;
lut[43] = 111;
lut[44] = 112;
lut[45] = 113;
lut[46] = 115;
lut[47] = 116;
lut[48] = 117;
lut[49] = 118;
lut[50] = 120;
lut[51] = 121;
lut[52] = 122;
lut[53] = 122;
lut[54] = 123;
lut[55] = 124;
lut[56] = 125;
lut[57] = 125;
lut[58] = 126;
lut[59] = 126;
lut[60] = 126;
lut[61] = 127;
lut[62] = 127;
lut[63] = 127;
lut[64] = 127;
lut[65] = 127;
lut[66] = 127;
lut[67] = 127;
lut[68] = 126;
lut[69] = 126;
lut[70] = 126;
lut[71] = 125;
lut[72] = 125;
lut[73] = 124;
lut[74] = 123;
lut[75] = 122;
lut[76] = 122;
lut[77] = 121;
lut[78] = 120;
lut[79] = 118;
lut[80] = 117;
lut[81] = 116;
lut[82] = 115;
lut[83] = 113;
lut[84] = 112;
lut[85] = 111;
lut[86] = 109;
lut[87] = 107;
lut[88] = 106;
lut[89] = 104;
lut[90] = 102;
lut[91] = 100;
lut[92] = 98;
lut[93] = 96;
lut[94] = 94;
lut[95] = 92;
lut[96] = 90;
lut[97] = 88;
lut[98] = 85;
lut[99] = 83;
lut[100] = 81;
lut[101] = 78;
lut[102] = 76;
lut[103] = 73;
lut[104] = 71;
lut[105] = 68;
lut[106] = 65;
lut[107] = 63;
lut[108] = 60;
lut[109] = 57;
lut[110] = 54;
lut[111] = 51;
lut[112] = 49;
lut[113] = 46;
lut[114] = 43;
lut[115] = 40;
lut[116] = 37;
lut[117] = 34;
lut[118] = 31;
lut[119] = 28;
lut[120] = 25;
lut[121] = 22;
lut[122] = 19;
lut[123] = 16;
lut[124] = 12;
lut[125] = 9;
lut[126] = 6;
lut[127] = 3;
lut[128] = 0;
lut[129] = -3;
lut[130] = -6;
lut[131] = -9;
lut[132] = -12;
lut[133] = -16;
lut[134] = -19;
lut[135] = -22;
lut[136] = -25;
lut[137] = -28;
lut[138] = -31;
lut[139] = -34;
lut[140] = -37;
lut[141] = -40;
lut[142] = -43;
lut[143] = -46;
lut[144] = -49;
lut[145] = -51;
lut[146] = -54;
lut[147] = -57;
lut[148] = -60;
lut[149] = -63;
lut[150] = -65;
lut[151] = -68;
lut[152] = -71;
lut[153] = -73;
lut[154] = -76;
lut[155] = -78;
lut[156] = -81;
lut[157] = -83;
lut[158] = -85;
lut[159] = -88;
lut[160] = -90;
lut[161] = -92;
lut[162] = -94;
lut[163] = -96;
lut[164] = -98;
lut[165] = -100;
lut[166] = -102;
lut[167] = -104;
lut[168] = -106;
lut[169] = -107;
lut[170] = -109;
lut[171] = -111;
lut[172] = -112;
lut[173] = -113;
lut[174] = -115;
lut[175] = -116;
lut[176] = -117;
lut[177] = -118;
lut[178] = -120;
lut[179] = -121;
lut[180] = -122;
lut[181] = -122;
lut[182] = -123;
lut[183] = -124;
lut[184] = -125;
lut[185] = -125;
lut[186] = -126;
lut[187] = -126;
lut[188] = -126;
lut[189] = -127;
lut[190] = -127;
lut[191] = -127;
lut[192] = -127;
lut[193] = -127;
lut[194] = -127;
lut[195] = -127;
lut[196] = -126;
lut[197] = -126;
lut[198] = -126;
lut[199] = -125;
lut[200] = -125;
lut[201] = -124;
lut[202] = -123;
lut[203] = -122;
lut[204] = -122;
lut[205] = -121;
lut[206] = -120;
lut[207] = -118;
lut[208] = -117;
lut[209] = -116;
lut[210] = -115;
lut[211] = -113;
lut[212] = -112;
lut[213] = -111;
lut[214] = -109;
lut[215] = -107;
lut[216] = -106;
lut[217] = -104;
lut[218] = -102;
lut[219] = -100;
lut[220] = -98;
lut[221] = -96;
lut[222] = -94;
lut[223] = -92;
lut[224] = -90;
lut[225] = -88;
lut[226] = -85;
lut[227] = -83;
lut[228] = -81;
lut[229] = -78;
lut[230] = -76;
lut[231] = -73;
lut[232] = -71;
lut[233] = -68;
lut[234] = -65;
lut[235] = -63;
lut[236] = -60;
lut[237] = -57;
lut[238] = -54;
lut[239] = -51;
lut[240] = -49;
lut[241] = -46;
lut[242] = -43;
lut[243] = -40;
lut[244] = -37;
lut[245] = -34;
lut[246] = -31;
lut[247] = -28;
lut[248] = -25;
lut[249] = -22;
lut[250] = -19;
lut[251] = -16;
lut[252] = -12;
lut[253] = -9;
lut[254] = -6;
lut[255] = -3;
     */
end

always @(posedge clk or posedge rst) begin
    if (rst) begin
        phase_acc <= phase;
        out <= 0;
        phase_increment <= 13;//freq_out*2^N/freq_clock, N-����������� lut(256=2^8)
    end else begin
        phase_acc <= phase_acc + phase_increment; 
        out <= lut[phase_acc[7:0]]; 
    end
end
endmodule